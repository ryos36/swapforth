//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.05
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9C
//Created Time: Tue Aug  9 16:53:52 2022

module Gowin_DPB (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [15:0] douta;
output [15:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [11:0] ada;
input [15:0] dina;
input [11:0] adb;
input [15:0] dinb;

wire [11:0] dpb_inst_0_douta_w;
wire [11:0] dpb_inst_0_doutb_w;
wire [11:0] dpb_inst_1_douta_w;
wire [11:0] dpb_inst_1_doutb_w;
wire [11:0] dpb_inst_2_douta_w;
wire [11:0] dpb_inst_2_doutb_w;
wire [11:0] dpb_inst_3_douta_w;
wire [11:0] dpb_inst_3_doutb_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[11:0],douta[3:0]}),
    .DOB({dpb_inst_0_doutb_w[11:0],doutb[3:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3:0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b0;
defparam dpb_inst_0.READ_MODE1 = 1'b0;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 4;
defparam dpb_inst_0.BIT_WIDTH_1 = 4;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'h6F31CF0E22A0E28F0C20F01610C3CC3E20F2C556F0D2CF1D2E5051564F1B2049;
defparam dpb_inst_0.INIT_RAM_01 = 256'h5A209814D4AC0007536630002F548F9103F00214936EFC1000314936ED00F3F3;
defparam dpb_inst_0.INIT_RAM_02 = 256'hD83016C74387C268222A8309377063A13FE941A981243546C0C2899DA22C9030;
defparam dpb_inst_0.INIT_RAM_03 = 256'h5CD03C0120D10440CDF10444F3F458D0B548F070424ACD07F3EC05242C03154C;
defparam dpb_inst_0.INIT_RAM_04 = 256'hF3F1FC8D31412EFF000000000310C1022401130CF837193C2DD4775F5CF07013;
defparam dpb_inst_0.INIT_RAM_05 = 256'h006F4F561F43C0F9300F4454AF514C06B9B014594EC03EF6E2001EF54DD33C10;
defparam dpb_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_07 = 256'h370B24C0557C7891C3D0371E237EE5540C9F1232FE62ABC171D4F50FEC000000;
defparam dpb_inst_0.INIT_RAM_08 = 256'h12301D798C00331301023A63030DEB26F1E36D9F13140F60C0047E74F3D10310;
defparam dpb_inst_0.INIT_RAM_09 = 256'h7C300004DD6ACD0503120313D1D7E7218D7B0B71A22F718F7777000D2D34CDD0;
defparam dpb_inst_0.INIT_RAM_0A = 256'h737C5873BCC55BC6075D55C6BB2121014733FFF432C4F303F03F1F303A311CD1;
defparam dpb_inst_0.INIT_RAM_0B = 256'h3D7730727F76821515DE74F7130337A01330A913C761031C061335471DE654DC;
defparam dpb_inst_0.INIT_RAM_0C = 256'h2263ED5311231171C1E6D6A6CC575D5121717046D5C6CC55113147C944CF023D;
defparam dpb_inst_0.INIT_RAM_0D = 256'h932364FA71F692251D31ACCC0080812176BF1D411B921252F6CDCD012CC0CC10;
defparam dpb_inst_0.INIT_RAM_0E = 256'h1BDE662BB1421C2CB300CC0F8E7153C2272D3169CFC5C9871922D2315411F0D3;
defparam dpb_inst_0.INIT_RAM_0F = 256'h64ED01EEDEE7E6C169019DA34A1ED031C1F495D96D0E31BDDE3E3CAC24C81C77;
defparam dpb_inst_0.INIT_RAM_10 = 256'h84FCE9553B03625B031851CDA9CFDE15BCCD7E3B30F130C7E54847F2EC7D6DD3;
defparam dpb_inst_0.INIT_RAM_11 = 256'hD8B4EBD655DB7B9F23C0484F0D61773DC03557FDC6F0D3F52E09E59B975B90BE;
defparam dpb_inst_0.INIT_RAM_12 = 256'hDC0BDFC51C91D34631D341F1C0D83AD0B0C1314DC8BD0F45C03121B4C0943BC0;
defparam dpb_inst_0.INIT_RAM_13 = 256'h222FE3AFF34F1EF16CF2ECA2EDEA1957CC0BD0FE638787781DDDD1280331D1E9;
defparam dpb_inst_0.INIT_RAM_14 = 256'h102FBDE25B722BD4550C0F38F93ED2644F024CD532C074AFC24F1EF12C45E6AF;
defparam dpb_inst_0.INIT_RAM_15 = 256'hD8F0372EFDE2D2000CD9C43613D2177966116829F225683D9285C52852CC558B;
defparam dpb_inst_0.INIT_RAM_16 = 256'hF8BCE0FCB0209E15977F405253AC4223252AE232092483208133F3725D0577FC;
defparam dpb_inst_0.INIT_RAM_17 = 256'h211CD619829891670053D6111D498B804A8DABC22084231284AC82CF061615F4;
defparam dpb_inst_0.INIT_RAM_18 = 256'h23C133D00AD27608D55011791967031109F183C0F037090079EF74536AC91030;
defparam dpb_inst_0.INIT_RAM_19 = 256'h73F8E10000000F5B170479FB2735454A4DD9D7B47277251C68044B4B01CC956C;
defparam dpb_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000088324728F4E42C11DB72129EA19C32AC;
defparam dpb_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_1 (
    .DOA({dpb_inst_1_douta_w[11:0],douta[7:4]}),
    .DOB({dpb_inst_1_doutb_w[11:0],doutb[7:4]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7:4]})
);

defparam dpb_inst_1.READ_MODE0 = 1'b0;
defparam dpb_inst_1.READ_MODE1 = 1'b0;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 4;
defparam dpb_inst_1.BIT_WIDTH_1 = 4;
defparam dpb_inst_1.BLK_SEL_0 = 3'b000;
defparam dpb_inst_1.BLK_SEL_1 = 3'b000;
defparam dpb_inst_1.RESET_MODE = "SYNC";
defparam dpb_inst_1.INIT_RAM_00 = 256'h7830681306203058030581042030380303806602803018020000666008020069;
defparam dpb_inst_1.INIT_RAM_01 = 256'h0E40760760D8507660C200500360A85110F01617670884110151767073108460;
defparam dpb_inst_1.INIT_RAM_02 = 256'h1B000682767058970589702703A3A001009501950140760182600770070F7267;
defparam dpb_inst_1.INIT_RAM_03 = 256'h0E310BE20E91760D89E1760C80660B91670AB121770991126088067088076078;
defparam dpb_inst_1.INIT_RAM_04 = 256'hF0F4F4030022038F000000003001B1403101602881011600011F22660FBD2D67;
defparam dpb_inst_1.INIT_RAM_05 = 256'h042B760E0B70D0B60D0B770C0B660A0E57461567099076608210066063100B10;
defparam dpb_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_07 = 256'h02120E8006660CE090110216770B7660B0B216098CC85411D17660F8FB000000;
defparam dpb_inst_1.INIT_RAM_08 = 256'h640012233901000001030410304F1203213020B21760181E0107660F80111011;
defparam dpb_inst_1.INIT_RAM_09 = 256'h29066666660A81101017001011221266114D1D2120A840883333D003C60581F0;
defparam dpb_inst_1.INIT_RAM_0A = 256'hFE660EF0418CBC0EA2010C0EA82121B15200777B021F88188901180201041911;
defparam dpb_inst_1.INIT_RAM_0B = 256'h01425E6028F1D2101666088610300226100023188CC1000B1B100D9D1766073F;
defparam dpb_inst_1.INIT_RAM_0C = 256'h05E02130112011213137602E0102013121212D57600E0003111152660D8EF021;
defparam dpb_inst_1.INIT_RAM_0D = 256'h50802F5B215BE75662760A806F60B121215823E809404067608313E207B1B114;
defparam dpb_inst_1.INIT_RAM_0E = 256'h141BEBA4B15A12049000267603903E203903E02FF66007021E753C760D268E10;
defparam dpb_inst_1.INIT_RAM_0F = 256'hE4F3017B6660DEC0DE00C3D0400A3100B17766608307B7973FEBBA767760682F;
defparam dpb_inst_1.INIT_RAM_10 = 256'h60687660690E60590E660483F2E7E0019883010100F100B018770E8078230110;
defparam dpb_inst_1.INIT_RAM_11 = 256'h3098791760D923660BAC408813012281A87760931B7017609A0660896607F136;
defparam dpb_inst_1.INIT_RAM_12 = 256'h4A5916602831102B01102B21A030093131B1A184A191760080007473A0660E80;
defparam dpb_inst_1.INIT_RAM_13 = 256'h70F860E860E80D80D820C820B3C06660AA09176609B2D22D1111108B10811069;
defparam dpb_inst_1.INIT_RAM_14 = 256'h14069130692705976058560486039770387702970297701830180080087660F8;
defparam dpb_inst_1.INIT_RAM_15 = 256'h11660262E3D62000081E02021012125B1C70AB0737609B01B760807608866079;
defparam dpb_inst_1.INIT_RAM_16 = 256'h6058A0FB90B0B16660B897C200A8F80A628096281962800181008022E17E268E;
defparam dpb_inst_1.INIT_RAM_17 = 256'h2118F1170870F1EEE0006CF17DDDBAB540B30CABB1D92077607A5BC2611C7667;
defparam dpb_inst_1.INIT_RAM_18 = 256'h80010001001F23001031112712173011331100107201007027107766098F280C;
defparam dpb_inst_1.INIT_RAM_19 = 256'h707B710508050F6660C688668E04770951151E45272256667084EC5081066600;
defparam dpb_inst_1.INIT_RAM_1A = 256'h00000000000000000000000000000000B907E87CB76008B118291873917370D8;
defparam dpb_inst_1.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_2 (
    .DOA({dpb_inst_2_douta_w[11:0],douta[11:8]}),
    .DOB({dpb_inst_2_doutb_w[11:0],doutb[11:8]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[11:8]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[11:8]})
);

defparam dpb_inst_2.READ_MODE0 = 1'b0;
defparam dpb_inst_2.READ_MODE1 = 1'b0;
defparam dpb_inst_2.WRITE_MODE0 = 2'b00;
defparam dpb_inst_2.WRITE_MODE1 = 2'b00;
defparam dpb_inst_2.BIT_WIDTH_0 = 4;
defparam dpb_inst_2.BIT_WIDTH_1 = 4;
defparam dpb_inst_2.BLK_SEL_0 = 3'b000;
defparam dpb_inst_2.BLK_SEL_1 = 3'b000;
defparam dpb_inst_2.RESET_MODE = "SYNC";
defparam dpb_inst_2.INIT_RAM_00 = 256'h01010F1050000008000081E000E00670C020BC3070000C001006047E02001066;
defparam dpb_inst_2.INIT_RAM_01 = 256'h30000000950D00009B003D00009B010013F9100068201001A100068C00101019;
defparam dpb_inst_2.INIT_RAM_02 = 256'hB040010155551000E1002E102000080030000000000004C10002100000300051;
defparam dpb_inst_2.INIT_RAM_03 = 256'h21012000B1110521000005F111022111034101110FD11B11421600541005C610;
defparam dpb_inst_2.INIT_RAM_04 = 256'h0301000130003230999999991301000321688D2001118ED21BB0112621001007;
defparam dpb_inst_2.INIT_RAM_05 = 256'h0DD082620084200EE20051320003220010115100421204522112045320B430B6;
defparam dpb_inst_2.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_07 = 256'h211043A904E9131012B1C10794F31028300003131110110010132723F0000000;
defparam dpb_inst_2.INIT_RAM_08 = 256'h1280B21221A1230801AA4404D44120D40043420000244C0001651543CFB112B1;
defparam dpb_inst_2.INIT_RAM_09 = 256'h11122220FF540B101CB26FB4B02121222B2111150D412A41222200002A54AB10;
defparam dpb_inst_2.INIT_RAM_0A = 256'h11E9141210002000210B0000221B1025112022227100521212305230F0C001B1;
defparam dpb_inst_2.INIT_RAM_0B = 256'h2B212011112021130225E5F10C0C3101023100020210A3001200022201493502;
defparam dpb_inst_2.INIT_RAM_0C = 256'h26013B12B112B1103005F36003010B111B351015F36003011B35110C6502112B;
defparam dpb_inst_2.INIT_RAM_0D = 256'h3C1C003611361130DE52060031330B11103F0021C63333035360000026010000;
defparam dpb_inst_2.INIT_RAM_0E = 256'h21B20331351300373409059D3730110373001C7024C17371111302520601C0B1;
defparam dpb_inst_2.INIT_RAM_0F = 256'h3020301251FA733A730B702003D70140001514D9703133310212337015937011;
defparam dpb_inst_2.INIT_RAM_10 = 256'h54891E728301098301451800240134B83000441436F05004410957C010103BB1;
defparam dpb_inst_2.INIT_RAM_11 = 256'h033113B51C8314404838031C1031111B315232800219BE54830C4583E1180140;
defparam dpb_inst_2.INIT_RAM_12 = 256'h4393B0FB9001B204F1B204013803140141004014393B0FC970204444394FF870;
defparam dpb_inst_2.INIT_RAM_13 = 256'h0F934195289CD92B99029A029020CD349383B0FC590101102BBBBA90121BB994;
defparam dpb_inst_2.INIT_RAM_14 = 256'hB02A3B02A310EAE804AD009A00EA105FA10F4A004A1013AF05A8CA7DA6026994;
defparam dpb_inst_2.INIT_RAM_15 = 256'hB255015020A5010000B1003017B111500237A00004F1A02B0313A0B13AA3C3A3;
defparam dpb_inst_2.INIT_RAM_16 = 256'h30B036F5365652C24CA15501015505055050550505505201517037014B541130;
defparam dpb_inst_2.INIT_RAM_17 = 256'h12005000000050055A02125035550505030030355155113013B37550500230E0;
defparam dpb_inst_2.INIT_RAM_18 = 256'h0006470170B51670B011B21006016FB16000016700167000100610031B050030;
defparam dpb_inst_2.INIT_RAM_19 = 256'h616060D006D06FC334C600000516091C3BB3B5631111304515C020360030C62C;
defparam dpb_inst_2.INIT_RAM_1A = 256'h000000000000000000000000000000000610406C0099D000B616E0000E000EC0;
defparam dpb_inst_2.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DPB dpb_inst_3 (
    .DOA({dpb_inst_3_douta_w[11:0],douta[15:12]}),
    .DOB({dpb_inst_3_doutb_w[11:0],doutb[15:12]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[15:12]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[15:12]})
);

defparam dpb_inst_3.READ_MODE0 = 1'b0;
defparam dpb_inst_3.READ_MODE1 = 1'b0;
defparam dpb_inst_3.WRITE_MODE0 = 2'b00;
defparam dpb_inst_3.WRITE_MODE1 = 2'b00;
defparam dpb_inst_3.BIT_WIDTH_0 = 4;
defparam dpb_inst_3.BIT_WIDTH_1 = 4;
defparam dpb_inst_3.BLK_SEL_0 = 3'b000;
defparam dpb_inst_3.BLK_SEL_1 = 3'b000;
defparam dpb_inst_3.RESET_MODE = "SYNC";
defparam dpb_inst_3.INIT_RAM_00 = 256'h0662066070080306803066300833066030682660680306803006076606803044;
defparam dpb_inst_3.INIT_RAM_01 = 256'h70092480660669247600666A8076060466F66260667060466626066600686626;
defparam dpb_inst_3.INIT_RAM_02 = 256'h606A406667660040200432006808268668448644860806606806004880600866;
defparam dpb_inst_3.INIT_RAM_03 = 256'h3006644020660730662607306677306606700666062066667706807706866606;
defparam dpb_inst_3.INIT_RAM_04 = 256'h8680848268606068666666662686460600667606606266600664667730046477;
defparam dpb_inst_3.INIT_RAM_05 = 256'h0004676004670046300466700407600004426407706606760066877600666466;
defparam dpb_inst_3.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_07 = 256'h66606066466660086666666667201076002467606044444626577706F4000000;
defparam dpb_inst_3.INIT_RAM_08 = 256'h5268646446666686866260063600406006670024606606444666666066666666;
defparam dpb_inst_3.INIT_RAM_09 = 256'h6664444062706664666266666646464406446466060642064444488482706648;
defparam dpb_inst_3.INIT_RAM_0A = 256'h4466600644600464064640642446462646684442644464646268666868686666;
defparam dpb_inst_3.INIT_RAM_0B = 256'h6646445466244462676730656686684866684864604066846466624265667008;
defparam dpb_inst_3.INIT_RAM_0C = 256'h3006064666466664260666006046464646266446660060446626460660604446;
defparam dpb_inst_3.INIT_RAM_0D = 256'h4656444866484540666770660426464660468085500808067700444030064460;
defparam dpb_inst_3.INIT_RAM_0E = 256'h646040442644607006C606666008440600844200876600866454486770056466;
defparam dpb_inst_3.INIT_RAM_0F = 256'h0484865466630043008500884850066846566666008544454844048066670664;
defparam dpb_inst_3.INIT_RAM_10 = 256'h6706566600A4060084666060824544300E64406266966C442506606856648666;
defparam dpb_inst_3.INIT_RAM_11 = 256'h084554E66600E4406008485664866656056767004456636600A6770066600640;
defparam dpb_inst_3.INIT_RAM_12 = 256'h4484E76206066660666662460848604646462654484E06606868044448463068;
defparam dpb_inst_3.INIT_RAM_13 = 256'h060666067706206206030603008866660084E066700646646666660066566600;
defparam dpb_inst_3.INIT_RAM_14 = 256'hE0700E0700E03066760664606760606606066067606067060706306306077606;
defparam dpb_inst_3.INIT_RAM_15 = 256'h6454664844848488066446646664660244420084876600660766002660676600;
defparam dpb_inst_3.INIT_RAM_16 = 256'h770606F04E462467760640044624408248082480824806864668668406446564;
defparam dpb_inst_3.INIT_RAM_17 = 256'h4646246484482600464654264000000408408440462406406600842444644067;
defparam dpb_inst_3.INIT_RAM_18 = 256'h0662668668646268644666646245266624868626886268486482507660624868;
defparam dpb_inst_3.INIT_RAM_19 = 256'h06042666C2666F67770044884464067006646444656640776600844486806670;
defparam dpb_inst_3.INIT_RAM_1A = 256'h0000000000000000000000000000000005644440406606066462644846480206;
defparam dpb_inst_3.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam dpb_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //Gowin_DPB
