`define UART_MASTER_SYSCLK 6.3e+07
`define UART_BAUD_RATE 115200
`define EBR_BASED
